typedef struct packed {
    logic [6:0] some_field;
} my_struct_t;

