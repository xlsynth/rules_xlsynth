localparam bit unsigned [31:0] Mol = 32'h0000002a;

typedef struct packed {
    logic [6:0] some_field;
} my_struct_t;

