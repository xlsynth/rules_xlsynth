module __main__main(
  input wire clk,
  output wire [31:0] out
);
  // ===== Pipe stage 0:
  assign out = 32'h0000_0040;
endmodule

